** Profile: "SCHEMATIC1-MCU_Power_Button"  [ c:\users\student\desktop\wcsa_sdp_2022\wcsa_orcad\pspice\mcu_powerbutton_simulation\mcu_power_button-pspicefiles\schematic1\mcu_power_button.sim ] 

** Creating circuit file "MCU_Power_Button.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../mcu_power_button-pspicefiles/mcu_power_button.lib" 
* From [PSPICE NETLIST] section of C:\Users\student\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\17.4.0\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 60 0 1m 
.OPTIONS ADVCONV
.PROBE64 V(*) I(*) W(*) D(*) NOISE(*) 
.INC "..\SCHEMATIC1.net" 


.END
