** Profile: "SCHEMATIC1-MCU_Power_Button"  [ C:\USERS\STUDENT\ORCAD_PCB\WCSA_ORCAD\MCU_POWERBUTTON_SIMULATION\mcu_power_button-pspicefiles\schematic1\mcu_power_button.sim ] 

** Creating circuit file "MCU_Power_Button.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../mcu_power_button-pspicefiles/mcu_power_button.lib" 
* From [PSPICE NETLIST] section of C:\Users\student\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\17.4.0\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 60 0 1m 
.OPTIONS ADVCONV
.PROBE64 V(*) I(*) W(*) D(*) NOISE(*) 
.INC "..\SCHEMATIC1.net" 


.END
