** Profile: "SCHEMATIC1-PowerBlock_Sim"  [ C:\Users\student\Desktop\WCSA_SDP_2022\WCSA_OrCAD\PSPICE\PowerSystem_Simulations\powersystem_simulations-pspicefiles\schematic1\powerblock_sim.sim ] 

** Creating circuit file "PowerBlock_Sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../powersystem_simulations-pspicefiles/powersystem_simulations.lib" 
.LIB "../../../powersystem_simulations-pspicefiles/schematic1/powerblock_sim/sllm359/mc33063a-q1_pspice_trans/mc33063a-q1_trans.lib"
+ "" 
* From [PSPICE NETLIST] section of C:\Users\student\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\17.4.0\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN 1e-03 6 0 50m 
.OPTIONS ADVCONV
.PROBE N([N87447])
.PROBE N([N37893])
.PROBE N([N44923])
.PROBE N([N87291])
.INC "..\SCHEMATIC1.net" 


.END
