** Profile: "SCHEMATIC1-PowerBlock_Sim"  [ C:\Users\student\OrCAD_PCB\WCSA_OrCAD\PowerSystem_Simulations\powersystem_simulations-pspicefiles\schematic1\powerblock_sim.sim ] 

** Creating circuit file "PowerBlock_Sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../powersystem_simulations-pspicefiles/powersystem_simulations.lib" 
.LIB "../../../powersystem_simulations-pspicefiles/schematic1/powerblock_sim/sllm359/mc33063a-q1_pspice_trans/mc33063a-q1_trans.lib"
+ "" 
* From [PSPICE NETLIST] section of C:\Users\student\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\17.4.0\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN 1e-03 500m 0 50m 
.OPTIONS ADVCONV
.PROBE64 N([N35320])
.PROBE64 N([N35162])
.PROBE64 N([N35460])
.PROBE64 N([N44923])
.INC "..\SCHEMATIC1.net" 


.END
